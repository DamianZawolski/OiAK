module mul3x3_17 (input a1,
                a2,
                a3,
                b1,
                b2,
                b3,
                output r1,
                r2,
                r3,
                r4,
                r5,
                r6);

    wire [1:6] p;
    assign p = {a1,a2,a3}*{b1,b2,b3};

    assign r1 = (!p[1]&p[2]&!p[4]&!p[5]&!p[6]) | (!p[1]&!p[2]&!p[3]&!p[4]&p[5]&!p[6]) | (
    p[1]&!p[2]&!p[3]&p[4]&p[5]&!p[6]) | (!p[1]&p[2]&!p[3]&!p[4]&p[5]&p[6]) | (
    !p[1]&p[2]&p[4]&p[5]&!p[6]) | (!p[1]&!p[2]&p[3]&!p[4]&!p[5]&!p[6]) | (
    p[1]&!p[2]&p[3]&p[4]&!p[5]&!p[6]) | (!p[1]&!p[2]&p[4]&!p[5]&p[6]) | (
    p[1]&!p[2]&!p[4]&!p[5]&p[6]) | (!p[1]&p[3]&!p[4]&p[5]&p[6]);

    assign r2 = (!p[1]&p[2]&!p[3]&!p[4]&p[5]&!p[6]) | (p[1]&!p[2]&!p[3]&p[4]&!p[5]
    &p[6]) | (!p[1]&!p[2]&p[3]&!p[4]&p[5]&!p[6]) | (!p[1]&p[2]&p[3]&!p[4]
    &p[5]&!p[6]) | (!p[1]&p[2]&p[4]&!p[5]&p[6]) | (!p[1]&!p[2]&!p[3]&!p[4]
    &!p[5]&p[6]) | (!p[1]&!p[2]&p[4]&!p[5]&!p[6]) | (p[1]&!p[2]&!p[4]
    &!p[5]&!p[6]) | (p[1]&!p[2]&p[3]&p[4]&p[5]&!p[6]) | (!p[1]&!p[2]&p[4]
    &p[5]&p[6]) | (p[1]&!p[2]&!p[4]&p[5]&p[6]);

    assign r3 = (!p[1]&p[2]&!p[3]&!p[4]&p[5]&!p[6]) | (p[1]&!p[2]&p[3]&p[4]&!p[5]
    &p[6]) | (!p[1]&p[2]&!p[3]&!p[4]&p[5]&p[6]) | (!p[1]&p[2]&!p[3]&p[4]
    &!p[5]&!p[6]) | (!p[1]&p[2]&p[4]&p[5]&!p[6]) | (!p[1]&!p[2]&p[3]&!p[4]
    &!p[5]&!p[6]) | (p[1]&!p[2]&p[3]&p[4]&!p[5]&!p[6]) | (p[1]&!p[2]&p[3]
    &p[4]&p[5]&!p[6]) | (p[1]&!p[2]&!p[4]&p[5]&p[6]) | (!p[1]&p[2]&!p[3]
    &p[4]&p[6]) | (!p[2]&p[3]&!p[4]&p[5]&!p[6]) | (!p[1]&p[2]&p[4]&p[5]
    &p[6]) | (p[1]&!p[2]&!p[3]&!p[4]) | (!p[1]&!p[2]&p[3]&!p[4]&p[6]) | (
    !p[1]&!p[3]&p[4]&p[5]);

    assign r4 = (p[1]&!p[2]&p[3]&p[4]&!p[5]&p[6]) | (!p[1]&!p[2]&p[3]&!p[4]&p[5]
    &!p[6]) | (!p[1]&!p[2]&!p[3]&p[4]&!p[5]&!p[6]) | (!p[1]&!p[2]&!p[3]
    &p[4]&!p[5]&p[6]) | (!p[2]&!p[3]&!p[4]&p[5]&p[6]) | (p[1]&!p[2]&p[3]
    &p[4]&p[5]&!p[6]) | (p[1]&!p[2]&!p[4]&!p[5]&p[6]) | (!p[1]&p[2]&p[3]
    &p[4]&!p[5]) | (!p[1]&!p[2]&p[3]&p[5]&p[6]) | (p[1]&!p[2]&p[3]&!p[4]
    &!p[5]) | (!p[1]&p[2]&!p[3]&p[4]&p[6]) | (!p[1]&p[2]&!p[3]&!p[4]&!p[5]) | (
    !p[1]&p[3]&!p[4]&p[5]&p[6]) | (!p[1]&p[2]&!p[3]&p[4]&p[5]) | (p[1]
    &!p[2]&!p[3]&!p[4]&p[5]) | (p[1]&!p[2]&!p[3]&p[5]&p[6]) | (!p[1]&!p[2]
    &p[3]&!p[4]&p[6]);

    assign r5 = (p[1]&!p[2]&!p[3]&p[4]&!p[5]&p[6]) | (!p[1]&p[2]&p[3]&!p[4]&p[5]
    &!p[6]) | (!p[1]&!p[2]&!p[3]&!p[4]&p[5]&!p[6]) | (p[1]&!p[2]&!p[3]
    &p[4]&p[5]&!p[6]) | (!p[1]&!p[2]&p[3]&p[4]&p[5]&!p[6]) | (!p[1]&p[2]
    &!p[3]&p[4]&!p[5]&!p[6]) | (!p[1]&p[2]&!p[4]&!p[5]&p[6]) | (!p[2]
    &p[3]&!p[4]&p[5]&p[6]) | (!p[1]&!p[2]&p[3]&!p[4]&!p[5]&!p[6]) | (
    !p[1]&!p[2]&!p[3]&p[4]&!p[5]&p[6]) | (p[1]&!p[2]&!p[4]&!p[5]&!p[6]) | (
    p[1]&!p[2]&p[3]&p[4]&!p[5]&!p[6]) | (p[1]&!p[2]&p[3]&p[4]&p[5]&!p[6]) | (
    !p[1]&p[2]&p[3]&p[4]&!p[5]) | (p[1]&!p[2]&p[3]&!p[4]&!p[5]) | (!p[1]
    &p[2]&p[4]&p[5]&p[6]) | (p[1]&!p[2]&!p[3]&!p[4]&p[5]);

    assign r6 = (p[1]&!p[2]&!p[3]&!p[5]&!p[6]) | (!p[1]&p[2]&p[3]&!p[4]&p[5]&!p[6]) | (
    p[1]&!p[2]&p[3]&!p[5]&p[6]) | (p[1]&!p[2]&!p[3]&p[4]&p[5]&!p[6]) | (
    !p[1]&p[2]&!p[3]&!p[4]&p[5]&p[6]) | (!p[1]&!p[2]&p[3]&p[4]&p[5]&!p[6]) | (
    !p[1]&!p[2]&!p[3]&!p[4]&!p[5]&p[6]) | (!p[1]&p[2]&!p[3]&p[4]&!p[5]
    &!p[6]) | (!p[1]&!p[2]&!p[3]&p[4]&!p[5]&!p[6]) | (!p[1]&p[3]&p[4]
    &!p[5]&p[6]) | (!p[1]&!p[3]&p[4]&p[5]&p[6]) | (p[1]&!p[2]&p[3]&p[4]
    &!p[5]&!p[6]) | (!p[2]&p[3]&!p[4]&p[5]&!p[6]) | (!p[1]&p[2]&!p[3]
    &!p[4]&!p[5]) | (!p[1]&p[2]&!p[3]&p[4]&p[5]) | (p[1]&!p[2]&!p[3]&p[5]
    &p[6]);

endmodule